magic
tech sky130B
magscale 1 2
timestamp 1714698450
<< error_p >>
rect -125 1199 -67 1205
rect 67 1199 125 1205
rect -125 1165 -113 1199
rect 67 1165 79 1199
rect -125 1159 -67 1165
rect 67 1159 125 1165
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -125 -1165 -67 -1159
rect 67 -1165 125 -1159
rect -125 -1199 -113 -1165
rect 67 -1199 79 -1165
rect -125 -1205 -67 -1199
rect 67 -1205 125 -1199
<< nwell >>
rect -311 -1337 311 1337
<< pmos >>
rect -111 118 -81 1118
rect -15 118 15 1118
rect 81 118 111 1118
rect -111 -1118 -81 -118
rect -15 -1118 15 -118
rect 81 -1118 111 -118
<< pdiff >>
rect -173 1106 -111 1118
rect -173 130 -161 1106
rect -127 130 -111 1106
rect -173 118 -111 130
rect -81 1106 -15 1118
rect -81 130 -65 1106
rect -31 130 -15 1106
rect -81 118 -15 130
rect 15 1106 81 1118
rect 15 130 31 1106
rect 65 130 81 1106
rect 15 118 81 130
rect 111 1106 173 1118
rect 111 130 127 1106
rect 161 130 173 1106
rect 111 118 173 130
rect -173 -130 -111 -118
rect -173 -1106 -161 -130
rect -127 -1106 -111 -130
rect -173 -1118 -111 -1106
rect -81 -130 -15 -118
rect -81 -1106 -65 -130
rect -31 -1106 -15 -130
rect -81 -1118 -15 -1106
rect 15 -130 81 -118
rect 15 -1106 31 -130
rect 65 -1106 81 -130
rect 15 -1118 81 -1106
rect 111 -130 173 -118
rect 111 -1106 127 -130
rect 161 -1106 173 -130
rect 111 -1118 173 -1106
<< pdiffc >>
rect -161 130 -127 1106
rect -65 130 -31 1106
rect 31 130 65 1106
rect 127 130 161 1106
rect -161 -1106 -127 -130
rect -65 -1106 -31 -130
rect 31 -1106 65 -130
rect 127 -1106 161 -130
<< nsubdiff >>
rect -275 1267 -179 1301
rect 179 1267 275 1301
rect -275 -1267 -241 1267
rect 241 -1267 275 1267
rect -275 -1301 275 -1267
<< nsubdiffcont >>
rect -179 1267 179 1301
<< poly >>
rect -129 1199 -63 1215
rect -129 1165 -113 1199
rect -79 1165 -63 1199
rect -129 1149 -63 1165
rect 63 1199 129 1215
rect 63 1165 79 1199
rect 113 1165 129 1199
rect 63 1149 129 1165
rect -111 1118 -81 1149
rect -15 1118 15 1144
rect 81 1118 111 1149
rect -111 92 -81 118
rect -15 87 15 118
rect 81 92 111 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -111 -118 -81 -92
rect -15 -118 15 -87
rect 81 -118 111 -92
rect -111 -1149 -81 -1118
rect -15 -1144 15 -1118
rect 81 -1149 111 -1118
rect -129 -1165 -63 -1149
rect -129 -1199 -113 -1165
rect -79 -1199 -63 -1165
rect -129 -1215 -63 -1199
rect 63 -1165 129 -1149
rect 63 -1199 79 -1165
rect 113 -1199 129 -1165
rect 63 -1215 129 -1199
<< polycont >>
rect -113 1165 -79 1199
rect 79 1165 113 1199
rect -17 37 17 71
rect -17 -71 17 -37
rect -113 -1199 -79 -1165
rect 79 -1199 113 -1165
<< locali >>
rect -195 1267 -179 1301
rect 179 1267 195 1301
rect -129 1165 -113 1199
rect -79 1165 -63 1199
rect 63 1165 79 1199
rect 113 1165 129 1199
rect -161 1106 -127 1122
rect -161 114 -127 130
rect -65 1106 -31 1122
rect -65 114 -31 130
rect 31 1106 65 1122
rect 31 114 65 130
rect 127 1106 161 1122
rect 127 114 161 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -161 -130 -127 -114
rect -161 -1122 -127 -1106
rect -65 -130 -31 -114
rect -65 -1122 -31 -1106
rect 31 -130 65 -114
rect 31 -1122 65 -1106
rect 127 -130 161 -114
rect 127 -1122 161 -1106
rect -129 -1199 -113 -1165
rect -79 -1199 -63 -1165
rect 63 -1199 79 -1165
rect 113 -1199 129 -1165
<< viali >>
rect -113 1165 -79 1199
rect 79 1165 113 1199
rect -161 179 -127 1057
rect -65 325 -31 911
rect 31 179 65 1057
rect 127 325 161 911
rect -17 37 17 71
rect -17 -71 17 -37
rect -161 -1057 -127 -179
rect -65 -911 -31 -325
rect 31 -1057 65 -179
rect 127 -911 161 -325
rect -113 -1199 -79 -1165
rect 79 -1199 113 -1165
<< metal1 >>
rect -125 1199 -67 1205
rect -125 1165 -113 1199
rect -79 1165 -67 1199
rect -125 1159 -67 1165
rect 67 1199 125 1205
rect 67 1165 79 1199
rect 113 1165 125 1199
rect 67 1159 125 1165
rect -167 1057 -121 1069
rect -167 179 -161 1057
rect -127 179 -121 1057
rect 25 1057 71 1069
rect -71 911 -25 923
rect -71 325 -65 911
rect -31 325 -25 911
rect -71 313 -25 325
rect -167 167 -121 179
rect 25 179 31 1057
rect 65 179 71 1057
rect 121 911 167 923
rect 121 325 127 911
rect 161 325 167 911
rect 121 313 167 325
rect 25 167 71 179
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -167 -179 -121 -167
rect -167 -1057 -161 -179
rect -127 -1057 -121 -179
rect 25 -179 71 -167
rect -71 -325 -25 -313
rect -71 -911 -65 -325
rect -31 -911 -25 -325
rect -71 -923 -25 -911
rect -167 -1069 -121 -1057
rect 25 -1057 31 -179
rect 65 -1057 71 -179
rect 121 -325 167 -313
rect 121 -911 127 -325
rect 161 -911 167 -325
rect 121 -923 167 -911
rect 25 -1069 71 -1057
rect -125 -1165 -67 -1159
rect -125 -1199 -113 -1165
rect -79 -1199 -67 -1165
rect -125 -1205 -67 -1199
rect 67 -1165 125 -1159
rect 67 -1199 79 -1165
rect 113 -1199 125 -1165
rect 67 -1205 125 -1199
<< properties >>
string FIXED_BBOX -258 -1284 258 1284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.15 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 90 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
