magic
tech sky130A
magscale 1 2
timestamp 1755204904
<< metal3 >>
rect -3216 1012 3216 1040
rect -3216 -1012 3132 1012
rect 3196 -1012 3216 1012
rect -3216 -1040 3216 -1012
<< via3 >>
rect 3132 -1012 3196 1012
<< mimcap >>
rect -3176 960 2824 1000
rect -3176 -960 -3136 960
rect 2784 -960 2824 960
rect -3176 -1000 2824 -960
<< mimcapcontact >>
rect -3136 -960 2784 960
<< metal4 >>
rect 3116 1012 3212 1028
rect -3137 960 2785 961
rect -3137 -960 -3136 960
rect 2784 -960 2785 960
rect -3137 -961 2785 -960
rect 3116 -1012 3132 1012
rect 3196 -1012 3212 1012
rect 3116 -1028 3212 -1012
<< labels >>
rlabel via3 3164 0 3164 0 0 C2
port 1 nsew
rlabel mimcapcontact -176 0 -176 0 0 C1
port 2 nsew
<< properties >>
string FIXED_BBOX -3216 -1040 2864 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 10 val 615.2 carea 2.00 cperi 0.19 class capacitor nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
