magic
tech sky130A
magscale 1 2
timestamp 1755201682
<< error_p >>
rect -29 -1511 29 -1505
rect -29 -1545 -17 -1511
rect -29 -1551 29 -1545
<< nwell >>
rect -211 -1684 211 1684
<< pmos >>
rect -15 -1464 15 1536
<< pdiff >>
rect -73 1524 -15 1536
rect -73 -1452 -61 1524
rect -27 -1452 -15 1524
rect -73 -1464 -15 -1452
rect 15 1524 73 1536
rect 15 -1452 27 1524
rect 61 -1452 73 1524
rect 15 -1464 73 -1452
<< pdiffc >>
rect -61 -1452 -27 1524
rect 27 -1452 61 1524
<< nsubdiff >>
rect -175 1614 -79 1648
rect 79 1614 175 1648
rect -175 -1614 -141 1614
rect 141 -1614 175 1614
rect -175 -1648 175 -1614
<< nsubdiffcont >>
rect -79 1614 79 1648
<< poly >>
rect -15 1536 15 1562
rect -15 -1495 15 -1464
rect -33 -1511 33 -1495
rect -33 -1545 -17 -1511
rect 17 -1545 33 -1511
rect -33 -1561 33 -1545
<< polycont >>
rect -17 -1545 17 -1511
<< locali >>
rect -95 1614 -79 1648
rect 79 1614 95 1648
rect -61 1524 -27 1540
rect -61 -1468 -27 -1452
rect 27 1524 61 1540
rect 27 -1468 61 -1452
rect -33 -1545 -17 -1511
rect 17 -1545 33 -1511
<< viali >>
rect -61 -1452 -27 1524
rect 27 -1006 61 1078
rect -17 -1545 17 -1511
<< metal1 >>
rect -67 1524 -21 1536
rect -67 -1452 -61 1524
rect -27 -1452 -21 1524
rect 21 1078 67 1090
rect 21 -1006 27 1078
rect 61 -1006 67 1078
rect 21 -1018 67 -1006
rect -67 -1464 -21 -1452
rect -29 -1511 29 -1505
rect -29 -1545 -17 -1511
rect 17 -1545 29 -1511
rect -29 -1551 29 -1545
<< labels >>
rlabel nsubdiff 0 -1631 0 -1631 0 B
port 1 nsew
rlabel pdiffc -44 36 -44 36 0 D
port 2 nsew
rlabel pdiffc 44 36 44 36 0 S
port 3 nsew
rlabel polycont 0 -1528 0 -1528 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -1631 158 1631
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 15 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
