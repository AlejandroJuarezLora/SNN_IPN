magic
tech sky130B
magscale 1 2
timestamp 1698529635
<< error_p >>
rect -29 249 29 255
rect -29 215 -17 249
rect -29 209 29 215
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect -29 -147 29 -141
rect -29 -463 29 -457
rect -29 -497 -17 -463
rect -29 -503 29 -497
<< pwell >>
rect -211 -635 211 635
<< nmos >>
rect -15 287 15 487
rect -15 -69 15 131
rect -15 -425 15 -225
<< ndiff >>
rect -73 475 -15 487
rect -73 299 -61 475
rect -27 299 -15 475
rect -73 287 -15 299
rect 15 475 73 487
rect 15 299 27 475
rect 61 299 73 475
rect 15 287 73 299
rect -73 119 -15 131
rect -73 -57 -61 119
rect -27 -57 -15 119
rect -73 -69 -15 -57
rect 15 119 73 131
rect 15 -57 27 119
rect 61 -57 73 119
rect 15 -69 73 -57
rect -73 -237 -15 -225
rect -73 -413 -61 -237
rect -27 -413 -15 -237
rect -73 -425 -15 -413
rect 15 -237 73 -225
rect 15 -413 27 -237
rect 61 -413 73 -237
rect 15 -425 73 -413
<< ndiffc >>
rect -61 299 -27 475
rect 27 299 61 475
rect -61 -57 -27 119
rect 27 -57 61 119
rect -61 -413 -27 -237
rect 27 -413 61 -237
<< psubdiff >>
rect -175 565 175 599
rect -175 -565 -141 565
rect 141 -565 175 565
rect -175 -599 -79 -565
rect 79 -599 175 -565
<< psubdiffcont >>
rect -79 -599 79 -565
<< poly >>
rect -15 487 15 513
rect -15 265 15 287
rect -33 249 33 265
rect -33 215 -17 249
rect 17 215 33 249
rect -33 199 33 215
rect -15 131 15 157
rect -15 -91 15 -69
rect -33 -107 33 -91
rect -33 -141 -17 -107
rect 17 -141 33 -107
rect -33 -157 33 -141
rect -15 -225 15 -199
rect -15 -447 15 -425
rect -33 -463 33 -447
rect -33 -497 -17 -463
rect 17 -497 33 -463
rect -33 -513 33 -497
<< polycont >>
rect -17 215 17 249
rect -17 -141 17 -107
rect -17 -497 17 -463
<< locali >>
rect -61 475 -27 491
rect -61 283 -27 299
rect 27 475 61 491
rect 27 283 61 299
rect -33 215 -17 249
rect 17 215 33 249
rect -61 119 -27 135
rect -61 -73 -27 -57
rect 27 119 61 135
rect 27 -73 61 -57
rect -33 -141 -17 -107
rect 17 -141 33 -107
rect -61 -237 -27 -221
rect -61 -429 -27 -413
rect 27 -237 61 -221
rect 27 -429 61 -413
rect -33 -497 -17 -463
rect 17 -497 33 -463
rect -95 -599 -79 -565
rect 79 -599 95 -565
<< viali >>
rect -61 299 -27 475
rect 27 334 61 440
rect -17 215 17 249
rect -61 -57 -27 119
rect 27 -22 61 84
rect -17 -141 17 -107
rect -61 -413 -27 -237
rect 27 -378 61 -272
rect -17 -497 17 -463
<< metal1 >>
rect -67 475 -21 487
rect -67 299 -61 475
rect -27 299 -21 475
rect 21 440 67 452
rect 21 334 27 440
rect 61 334 67 440
rect 21 322 67 334
rect -67 287 -21 299
rect -29 249 29 255
rect -29 215 -17 249
rect 17 215 29 249
rect -29 209 29 215
rect -67 119 -21 131
rect -67 -57 -61 119
rect -27 -57 -21 119
rect 21 84 67 96
rect 21 -22 27 84
rect 61 -22 67 84
rect 21 -34 67 -22
rect -67 -69 -21 -57
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect 17 -141 29 -107
rect -29 -147 29 -141
rect -67 -237 -21 -225
rect -67 -413 -61 -237
rect -27 -413 -21 -237
rect 21 -272 67 -260
rect 21 -378 27 -272
rect 61 -378 67 -272
rect 21 -390 67 -378
rect -67 -425 -21 -413
rect -29 -463 29 -457
rect -29 -497 -17 -463
rect 17 -497 29 -463
rect -29 -503 29 -497
<< properties >>
string FIXED_BBOX -158 -582 158 582
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
