* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_pr_reram__reram_cell_london TE BE
N1 TE BE sky130_fd_pr_reram__reram_cell_london_model
.ends sky130_fd_pr_reram__reram_cell_london



.model sky130_fd_pr_reram__reram_cell_london_model sky130_fd_pr_reram__reram_cell_london_va 

.control
pre_osdi /home/alex/pdk/sky130B/libs.tech/ngspice/sky130_fd_pr_reram__reram_cell_london.osdi
.endc

