magic
tech sky130B
magscale 1 2
timestamp 1714698238
<< error_p >>
rect -77 1699 -19 1705
rect -77 1665 -65 1699
rect -77 1659 -19 1665
rect 19 71 77 77
rect 19 37 31 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 19 -77 77 -71
rect -77 -1665 -19 -1659
rect -77 -1699 -65 -1665
rect -77 -1705 -19 -1699
<< nwell >>
rect -263 -1837 263 1837
<< pmos >>
rect -63 118 -33 1618
rect 33 118 63 1618
rect -63 -1618 -33 -118
rect 33 -1618 63 -118
<< pdiff >>
rect -125 1606 -63 1618
rect -125 130 -113 1606
rect -79 130 -63 1606
rect -125 118 -63 130
rect -33 1606 33 1618
rect -33 130 -17 1606
rect 17 130 33 1606
rect -33 118 33 130
rect 63 1606 125 1618
rect 63 130 79 1606
rect 113 130 125 1606
rect 63 118 125 130
rect -125 -130 -63 -118
rect -125 -1606 -113 -130
rect -79 -1606 -63 -130
rect -125 -1618 -63 -1606
rect -33 -130 33 -118
rect -33 -1606 -17 -130
rect 17 -1606 33 -130
rect -33 -1618 33 -1606
rect 63 -130 125 -118
rect 63 -1606 79 -130
rect 113 -1606 125 -130
rect 63 -1618 125 -1606
<< pdiffc >>
rect -113 130 -79 1606
rect -17 130 17 1606
rect 79 130 113 1606
rect -113 -1606 -79 -130
rect -17 -1606 17 -130
rect 79 -1606 113 -130
<< nsubdiff >>
rect -227 1767 -131 1801
rect 131 1767 227 1801
rect -227 -1767 -193 1767
rect 193 -1767 227 1767
rect -227 -1801 227 -1767
<< nsubdiffcont >>
rect -131 1767 131 1801
<< poly >>
rect -81 1699 -15 1715
rect -81 1665 -65 1699
rect -31 1665 -15 1699
rect -81 1649 -15 1665
rect -63 1618 -33 1649
rect 33 1618 63 1644
rect -63 92 -33 118
rect 33 87 63 118
rect 15 71 81 87
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 15 -87 81 -71
rect -63 -118 -33 -92
rect 33 -118 63 -87
rect -63 -1649 -33 -1618
rect 33 -1644 63 -1618
rect -81 -1665 -15 -1649
rect -81 -1699 -65 -1665
rect -31 -1699 -15 -1665
rect -81 -1715 -15 -1699
<< polycont >>
rect -65 1665 -31 1699
rect 31 37 65 71
rect 31 -71 65 -37
rect -65 -1699 -31 -1665
<< locali >>
rect -147 1767 -131 1801
rect 131 1767 147 1801
rect -81 1665 -65 1699
rect -31 1665 -15 1699
rect -113 1606 -79 1622
rect -113 114 -79 130
rect -17 1606 17 1622
rect -17 114 17 130
rect 79 1606 113 1622
rect 79 114 113 130
rect 15 37 31 71
rect 65 37 81 71
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -113 -130 -79 -114
rect -113 -1622 -79 -1606
rect -17 -130 17 -114
rect -17 -1622 17 -1606
rect 79 -130 113 -114
rect 79 -1622 113 -1606
rect -81 -1699 -65 -1665
rect -31 -1699 -15 -1665
<< viali >>
rect -65 1665 -31 1699
rect -113 204 -79 1532
rect -17 425 17 1311
rect 79 204 113 1532
rect 31 37 65 71
rect 31 -71 65 -37
rect -113 -1532 -79 -204
rect -17 -1311 17 -425
rect 79 -1532 113 -204
rect -65 -1699 -31 -1665
<< metal1 >>
rect -77 1699 -19 1705
rect -77 1665 -65 1699
rect -31 1665 -19 1699
rect -77 1659 -19 1665
rect -119 1532 -73 1544
rect -119 204 -113 1532
rect -79 204 -73 1532
rect 73 1532 119 1544
rect -23 1311 23 1323
rect -23 425 -17 1311
rect 17 425 23 1311
rect -23 413 23 425
rect -119 192 -73 204
rect 73 204 79 1532
rect 113 204 119 1532
rect 73 192 119 204
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect -119 -204 -73 -192
rect -119 -1532 -113 -204
rect -79 -1532 -73 -204
rect 73 -204 119 -192
rect -23 -425 23 -413
rect -23 -1311 -17 -425
rect 17 -1311 23 -425
rect -23 -1323 23 -1311
rect -119 -1544 -73 -1532
rect 73 -1532 79 -204
rect 113 -1532 119 -204
rect 73 -1544 119 -1532
rect -77 -1665 -19 -1659
rect -77 -1699 -65 -1665
rect -31 -1699 -19 -1665
rect -77 -1705 -19 -1699
<< properties >>
string FIXED_BBOX -210 -1784 210 1784
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.5 l 0.15 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 90 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
