magic
tech sky130A
magscale 1 2
timestamp 1757008927
<< nwell >>
rect -311 -703 311 703
<< pmos >>
rect -111 -483 -81 517
rect -15 -483 15 517
rect 81 -483 111 517
<< pdiff >>
rect -173 505 -111 517
rect -173 -471 -161 505
rect -127 -471 -111 505
rect -173 -483 -111 -471
rect -81 505 -15 517
rect -81 -471 -65 505
rect -31 -471 -15 505
rect -81 -483 -15 -471
rect 15 505 81 517
rect 15 -471 31 505
rect 65 -471 81 505
rect 15 -483 81 -471
rect 111 505 173 517
rect 111 -471 127 505
rect 161 -471 173 505
rect 111 -483 173 -471
<< pdiffc >>
rect -161 -471 -127 505
rect -65 -471 -31 505
rect 31 -471 65 505
rect 127 -471 161 505
<< nsubdiff >>
rect -275 633 -179 667
rect 179 633 275 667
rect -275 -633 -241 633
rect 241 -633 275 633
rect -275 -667 275 -633
<< nsubdiffcont >>
rect -179 633 179 667
<< poly >>
rect -111 517 -81 543
rect -15 517 15 581
rect 81 517 111 543
rect -111 -514 -81 -483
rect -15 -509 15 -483
rect 81 -514 111 -483
rect -129 -530 -63 -514
rect -129 -564 -113 -530
rect -79 -564 -63 -530
rect -129 -580 -63 -564
rect 63 -530 129 -514
rect 63 -564 79 -530
rect 113 -564 129 -530
rect 63 -580 129 -564
<< polycont >>
rect -113 -564 -79 -530
rect 79 -564 113 -530
<< locali >>
rect -195 633 -179 667
rect 179 633 195 667
rect -161 505 -127 521
rect -161 -487 -127 -471
rect -65 505 -31 521
rect -65 -487 -31 -471
rect 31 505 65 521
rect 31 -487 65 -471
rect 127 505 161 521
rect 127 -487 161 -471
rect -129 -564 -113 -530
rect -79 -564 -63 -530
rect 63 -564 79 -530
rect 113 -564 129 -530
<< viali >>
rect -161 -471 -127 505
rect -65 -325 -31 359
rect 31 -471 65 505
rect 127 -325 161 359
rect -113 -564 -79 -530
rect 79 -564 113 -530
<< metal1 >>
rect -163 517 69 539
rect -167 505 71 517
rect -167 -471 -161 505
rect -127 491 31 505
rect -127 -471 -121 491
rect -71 359 -25 371
rect -71 -248 -65 359
rect -76 -254 -65 -248
rect -31 -248 -25 359
rect -31 -254 -24 -248
rect -76 -312 -65 -306
rect -71 -325 -65 -312
rect -31 -312 -24 -306
rect -31 -325 -25 -312
rect -71 -337 -25 -325
rect -167 -483 -121 -471
rect 25 -471 31 491
rect 65 -471 71 505
rect 121 359 167 371
rect 121 -254 127 359
rect 161 -248 167 359
rect 161 -254 177 -248
rect 121 -306 125 -254
rect 177 -298 187 -262
rect 121 -325 127 -306
rect 161 -312 177 -306
rect 161 -325 167 -312
rect 121 -337 167 -325
rect 25 -483 71 -471
rect -125 -530 -67 -524
rect 67 -530 125 -524
rect -125 -564 -113 -530
rect -79 -564 79 -530
rect 113 -564 125 -530
rect -125 -570 -67 -564
rect 67 -570 125 -564
<< via1 >>
rect -76 -306 -65 -254
rect -65 -306 -31 -254
rect -31 -306 -24 -254
rect 125 -306 127 -254
rect 127 -306 161 -254
rect 161 -306 177 -254
<< metal2 >>
rect -82 -306 -76 -254
rect -24 -262 -18 -254
rect 119 -262 125 -254
rect -24 -298 125 -262
rect -24 -306 -18 -298
rect 119 -306 125 -298
rect 177 -306 183 -254
<< labels >>
flabel metal1 s -143 20 -143 20 0 FreeSans 320 0 0 0 D
port 0 nsew
flabel metal1 s 146 32 146 32 0 FreeSans 320 0 0 0 S
port 1 nsew
flabel metal1 s 0 -546 0 -546 0 FreeSans 320 0 0 0 G
port 2 nsew
flabel locali s 6 650 6 650 0 FreeSans 320 0 0 0 B
port 3 nsew
<< end >>
