magic
tech sky130A
magscale 1 2
timestamp 1755201682
<< error_p >>
rect -29 -411 29 -405
rect -29 -445 -17 -411
rect -29 -451 29 -445
<< nwell >>
rect -211 -584 211 584
<< pmos >>
rect -15 -364 15 436
<< pdiff >>
rect -73 424 -15 436
rect -73 -352 -61 424
rect -27 -352 -15 424
rect -73 -364 -15 -352
rect 15 424 73 436
rect 15 -352 27 424
rect 61 -352 73 424
rect 15 -364 73 -352
<< pdiffc >>
rect -61 -352 -27 424
rect 27 -352 61 424
<< nsubdiff >>
rect -175 514 -79 548
rect 79 514 175 548
rect -175 -514 -141 514
rect 141 -514 175 514
rect -175 -548 175 -514
<< nsubdiffcont >>
rect -79 514 79 548
<< poly >>
rect -15 436 15 462
rect -15 -395 15 -364
rect -33 -411 33 -395
rect -33 -445 -17 -411
rect 17 -445 33 -411
rect -33 -461 33 -445
<< polycont >>
rect -17 -445 17 -411
<< locali >>
rect -95 514 -79 548
rect 79 514 95 548
rect -61 424 -27 440
rect -61 -368 -27 -352
rect 27 424 61 440
rect 27 -368 61 -352
rect -33 -445 -17 -411
rect 17 -445 33 -411
<< viali >>
rect -61 -352 -27 424
rect 27 -236 61 308
rect -17 -445 17 -411
<< metal1 >>
rect -67 424 -21 436
rect -67 -352 -61 424
rect -27 -352 -21 424
rect 21 308 67 320
rect 21 -236 27 308
rect 61 -236 67 308
rect 21 -248 67 -236
rect -67 -364 -21 -352
rect -29 -411 29 -405
rect -29 -445 -17 -411
rect 17 -445 29 -411
rect -29 -451 29 -445
<< labels >>
rlabel nsubdiff 0 -531 0 -531 0 B
port 1 nsew
rlabel pdiffc -44 36 -44 36 0 D
port 2 nsew
rlabel pdiffc 44 36 44 36 0 S
port 3 nsew
rlabel polycont 0 -428 0 -428 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -531 158 531
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
