magic
tech sky130A
magscale 1 2
timestamp 1755201682
<< nwell >>
rect -1196 -284 1196 284
<< pmos >>
rect -1000 -64 1000 136
<< pdiff >>
rect -1058 124 -1000 136
rect -1058 -52 -1046 124
rect -1012 -52 -1000 124
rect -1058 -64 -1000 -52
rect 1000 124 1058 136
rect 1000 -52 1012 124
rect 1046 -52 1058 124
rect 1000 -64 1058 -52
<< pdiffc >>
rect -1046 -52 -1012 124
rect 1012 -52 1046 124
<< nsubdiff >>
rect -1160 214 1160 248
rect -1160 -214 -1126 214
rect 1126 -214 1160 214
rect -1160 -248 -1064 -214
rect 1064 -248 1160 -214
<< nsubdiffcont >>
rect -1064 -248 1064 -214
<< poly >>
rect -1000 136 1000 162
rect -1000 -111 1000 -64
rect -1000 -145 -984 -111
rect 984 -145 1000 -111
rect -1000 -161 1000 -145
<< polycont >>
rect -984 -145 984 -111
<< locali >>
rect -1046 124 -1012 140
rect -1046 -68 -1012 -52
rect 1012 124 1046 140
rect 1012 -68 1046 -52
rect -1000 -145 -984 -111
rect 984 -145 1000 -111
rect -1080 -248 -1064 -214
rect 1064 -248 1080 -214
<< viali >>
rect -1046 -52 -1012 124
rect 1012 -26 1046 98
rect -984 -145 984 -111
<< metal1 >>
rect -1052 124 -1006 136
rect -1052 -52 -1046 124
rect -1012 -52 -1006 124
rect 1006 98 1052 110
rect 1006 -26 1012 98
rect 1046 -26 1052 98
rect 1006 -38 1052 -26
rect -1052 -64 -1006 -52
rect -996 -111 996 -105
rect -996 -145 -984 -111
rect 984 -145 996 -111
rect -996 -151 996 -145
<< labels >>
rlabel nsubdiffcont 0 -231 0 -231 0 B
port 1 nsew
rlabel pdiffc -1029 36 -1029 36 0 D
port 2 nsew
rlabel pdiffc 1029 36 1029 36 0 S
port 3 nsew
rlabel polycont 0 -128 0 -128 0 G
port 4 nsew
<< properties >>
string FIXED_BBOX -1143 -231 1143 231
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
