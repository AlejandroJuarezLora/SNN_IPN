magic
tech sky130B
magscale 1 2
timestamp 1714756698
<< error_p >>
rect -125 381 -67 387
rect 67 381 125 387
rect -125 347 -113 381
rect 67 347 79 381
rect -125 341 -67 347
rect 67 341 125 347
rect -221 -347 -163 -341
rect -29 -347 29 -341
rect 163 -347 221 -341
rect -221 -381 -209 -347
rect -29 -381 -17 -347
rect 163 -381 175 -347
rect -221 -387 -163 -381
rect -29 -387 29 -381
rect 163 -387 221 -381
<< nwell >>
rect -407 -519 407 519
<< pmos >>
rect -207 -300 -177 300
rect -111 -300 -81 300
rect -15 -300 15 300
rect 81 -300 111 300
rect 177 -300 207 300
<< pdiff >>
rect -269 288 -207 300
rect -269 -288 -257 288
rect -223 -288 -207 288
rect -269 -300 -207 -288
rect -177 288 -111 300
rect -177 -288 -161 288
rect -127 -288 -111 288
rect -177 -300 -111 -288
rect -81 288 -15 300
rect -81 -288 -65 288
rect -31 -288 -15 288
rect -81 -300 -15 -288
rect 15 288 81 300
rect 15 -288 31 288
rect 65 -288 81 288
rect 15 -300 81 -288
rect 111 288 177 300
rect 111 -288 127 288
rect 161 -288 177 288
rect 111 -300 177 -288
rect 207 288 269 300
rect 207 -288 223 288
rect 257 -288 269 288
rect 207 -300 269 -288
<< pdiffc >>
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
<< nsubdiff >>
rect -371 449 -275 483
rect 275 449 371 483
rect -371 -449 -337 449
rect 337 -449 371 449
rect -371 -483 371 -449
<< nsubdiffcont >>
rect -275 449 275 483
<< poly >>
rect -129 381 -63 397
rect -129 347 -113 381
rect -79 347 -63 381
rect -129 331 -63 347
rect 63 381 129 397
rect 63 347 79 381
rect 113 347 129 381
rect 63 331 129 347
rect -207 300 -177 326
rect -111 300 -81 331
rect -15 300 15 326
rect 81 300 111 331
rect 177 300 207 326
rect -207 -331 -177 -300
rect -111 -326 -81 -300
rect -15 -331 15 -300
rect 81 -326 111 -300
rect 177 -331 207 -300
rect -225 -347 -159 -331
rect -225 -381 -209 -347
rect -175 -381 -159 -347
rect -225 -397 -159 -381
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect 159 -347 225 -331
rect 159 -381 175 -347
rect 209 -381 225 -347
rect 159 -397 225 -381
<< polycont >>
rect -113 347 -79 381
rect 79 347 113 381
rect -209 -381 -175 -347
rect -17 -381 17 -347
rect 175 -381 209 -347
<< locali >>
rect -291 449 -275 483
rect 275 449 291 483
rect -129 347 -113 381
rect -79 347 -63 381
rect 63 347 79 381
rect 113 347 129 381
rect -257 288 -223 304
rect -257 -304 -223 -288
rect -161 288 -127 304
rect -161 -304 -127 -288
rect -65 288 -31 304
rect -65 -304 -31 -288
rect 31 288 65 304
rect 31 -304 65 -288
rect 127 288 161 304
rect 127 -304 161 -288
rect 223 288 257 304
rect 223 -304 257 -288
rect -225 -381 -209 -347
rect -175 -381 -159 -347
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect 159 -381 175 -347
rect 209 -381 225 -347
<< viali >>
rect -113 347 -79 381
rect 79 347 113 381
rect -257 -259 -223 259
rect -161 -173 -127 173
rect -65 -259 -31 259
rect 31 -173 65 173
rect 127 -259 161 259
rect 223 -173 257 173
rect -209 -381 -175 -347
rect -17 -381 17 -347
rect 175 -381 209 -347
<< metal1 >>
rect -125 381 -67 387
rect -125 347 -113 381
rect -79 347 -67 381
rect -125 341 -67 347
rect 67 381 125 387
rect 67 347 79 381
rect 113 347 125 381
rect 67 341 125 347
rect -263 259 -217 271
rect -263 -259 -257 259
rect -223 -259 -217 259
rect -71 259 -25 271
rect -167 173 -121 185
rect -167 -173 -161 173
rect -127 -173 -121 173
rect -167 -185 -121 -173
rect -263 -271 -217 -259
rect -71 -259 -65 259
rect -31 -259 -25 259
rect 121 259 167 271
rect 25 173 71 185
rect 25 -173 31 173
rect 65 -173 71 173
rect 25 -185 71 -173
rect -71 -271 -25 -259
rect 121 -259 127 259
rect 161 -259 167 259
rect 217 173 263 185
rect 217 -173 223 173
rect 257 -173 263 173
rect 217 -185 263 -173
rect 121 -271 167 -259
rect -221 -347 -163 -341
rect -221 -381 -209 -347
rect -175 -381 -163 -347
rect -221 -387 -163 -381
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect 163 -347 221 -341
rect 163 -381 175 -347
rect 209 -381 221 -347
rect 163 -387 221 -381
<< properties >>
string FIXED_BBOX -354 -466 354 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 90 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
