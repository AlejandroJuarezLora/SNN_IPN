magic
tech sky130B
magscale 1 2
timestamp 1715117223
<< nwell >>
rect -272 867 1804 1244
<< nsubdiff >>
rect 423 1175 1132 1209
<< locali >>
rect 389 1175 1135 1209
rect -152 906 111 940
rect 77 839 111 906
rect 389 839 423 1175
rect 1101 939 1135 1175
rect 1101 905 1303 939
rect 1337 905 1618 939
rect 1652 905 1677 939
rect 77 805 423 839
rect -135 -844 -101 -735
rect 1041 -844 1075 -717
rect 1355 -844 1389 -744
rect 1671 -844 1705 -748
rect -168 -878 1739 -844
<< viali >>
rect 1303 905 1337 939
rect 1618 905 1652 939
<< metal1 >>
rect 1530 1001 1764 1033
rect 1297 939 1343 951
rect 1297 905 1303 939
rect 1337 905 1343 939
rect 1297 893 1343 905
rect 1303 750 1337 893
rect 1530 786 1562 1001
rect 1612 939 1658 951
rect 1612 905 1618 939
rect 1652 905 1658 939
rect 1612 893 1658 905
rect 1618 743 1652 893
rect -48 586 4 592
rect -207 547 -82 581
rect -48 528 4 534
rect 265 586 317 592
rect 265 528 317 534
rect 72 425 228 459
rect 388 457 542 491
rect -376 348 -44 382
rect -376 -877 -342 348
rect 72 272 106 425
rect 388 375 422 457
rect 1171 439 1248 471
rect 1171 427 1217 439
rect 258 341 569 375
rect -242 238 106 272
rect -242 32 -209 238
rect -242 -27 -210 32
rect 383 -19 417 341
rect 1171 178 1203 427
rect 1250 344 1256 396
rect 1308 344 1314 396
rect 1555 333 1561 393
rect 1621 333 1627 393
rect 1732 273 1764 1001
rect 1731 241 2052 273
rect 1171 146 1967 178
rect 374 -25 426 -19
rect -242 -177 -203 -27
rect 1800 -54 1806 -2
rect 1858 -54 1864 -2
rect 374 -83 426 -77
rect -242 -183 -192 -177
rect -242 -216 -155 -183
rect -242 -223 -180 -216
rect -242 -285 -210 -223
rect 1935 -284 1967 146
rect -242 -286 101 -285
rect -242 -319 268 -286
rect -242 -323 -210 -319
rect 67 -320 268 -319
rect -264 -537 -258 -485
rect -206 -494 -200 -485
rect -206 -528 -40 -494
rect -206 -537 -200 -528
rect 67 -579 101 -320
rect 234 -496 268 -320
rect 1472 -316 1967 -284
rect 225 -529 1362 -496
rect 225 -530 393 -529
rect 464 -530 1362 -529
rect -47 -613 101 -579
rect 163 -651 169 -599
rect 221 -651 227 -599
rect 1266 -764 1301 -750
rect 1266 -792 1307 -764
rect 1472 -792 1504 -316
rect 1609 -529 1615 -477
rect 1667 -529 1673 -477
rect 1583 -765 1615 -729
rect 1577 -792 1623 -765
rect 1266 -808 1504 -792
rect 1267 -824 1504 -808
rect 1576 -793 1623 -792
rect 2020 -793 2052 241
rect 1576 -824 2052 -793
rect 1577 -825 2052 -824
rect 1577 -877 1623 -825
rect -376 -881 1623 -877
rect -376 -911 1622 -881
rect -376 -912 -342 -911
rect 1578 -916 1622 -911
<< via1 >>
rect -48 534 4 586
rect 265 534 317 586
rect 1256 344 1308 396
rect 1561 333 1621 393
rect 374 -77 426 -25
rect 1806 -54 1858 -2
rect -258 -537 -206 -485
rect 169 -651 221 -599
rect 1615 -529 1667 -477
<< metal2 >>
rect -54 534 -48 586
rect 4 577 10 586
rect 259 577 265 586
rect 4 543 265 577
rect 4 534 10 543
rect 259 534 265 543
rect 317 577 323 586
rect 317 543 1139 577
rect 317 534 323 543
rect 1105 173 1139 543
rect 1256 396 1308 402
rect 1561 393 1621 399
rect 1308 347 1362 393
rect 1256 338 1308 344
rect 1621 339 1983 387
rect 1561 327 1621 333
rect 1105 139 1849 173
rect 1815 4 1849 139
rect 1806 -2 1858 4
rect 368 -34 374 -25
rect 178 -68 374 -34
rect -258 -485 -206 -479
rect -258 -543 -206 -537
rect 178 -593 212 -68
rect 368 -77 374 -68
rect 426 -77 432 -25
rect 1806 -60 1858 -54
rect 1615 -477 1667 -471
rect 1935 -490 1983 339
rect 1667 -526 1983 -490
rect 1615 -535 1667 -529
rect 1935 -532 1983 -526
rect 169 -599 221 -593
rect 169 -657 221 -651
use M5  M5_0
timestamp 1715104367
transform -1 0 -73 0 1 -635
box -211 -279 211 279
use M5  M5_1
timestamp 1715104367
transform 1 0 1328 0 1 -635
box -211 -279 211 279
use M6  M6_0
timestamp 1715103727
transform -1 0 -62 0 1 591
box -211 -384 211 384
use M6  M6_1
timestamp 1715103727
transform 1 0 1591 0 1 591
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_GSRC26  sky130_fd_pr__nfet_01v8_GSRC26_0
timestamp 1715109623
transform 1 0 627 0 -1 -636
box -596 -241 601 279
use M5  sky130_fd_pr__nfet_01v8_NE5NAH_0
timestamp 1715104367
transform 1 0 1644 0 1 -635
box -211 -279 211 279
use M3  sky130_fd_pr__pfet_01v8_9RBQXV_0
timestamp 1715103490
transform 1 0 762 0 1 726
box -407 -519 407 519
use M1  sky130_fd_pr__pfet_01v8_AXGCW8_0
timestamp 1715102943
transform 1 0 803 0 1 -72
box -1196 -284 1196 284
use M2  sky130_fd_pr__pfet_01v8_HERV5D_0
timestamp 1715103109
transform 1 0 251 0 1 541
box -211 -334 211 334
use M6  sky130_fd_pr__pfet_01v8_MNLW5D_0
timestamp 1715103727
transform 1 0 1276 0 1 591
box -211 -384 211 384
<< labels >>
flabel locali s 468 1196 468 1196 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal2 379 557 379 557 0 FreeSans 480 0 0 0 vm
flabel metal1 -207 547 -82 581 0 FreeSans 480 0 0 0 Iext
port 1 nsew
flabel locali -168 -878 1739 -844 0 FreeSans 480 0 0 0 vss
port 2 nsew
flabel metal1 2008 251 2008 251 0 FreeSans 480 0 0 0 vout
port 5 nsew
flabel metal1 84 -372 84 -372 0 FreeSans 480 0 0 0 vg
flabel metal2 1316 347 1362 393 0 FreeSans 480 0 0 0 vb2
port 6 nsew
flabel via1 -233 -513 -233 -513 0 FreeSans 480 0 0 0 vb2
port 7 nsew
<< end >>
