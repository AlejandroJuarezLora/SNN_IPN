magic
tech sky130B
magscale 1 2
timestamp 1715103490
<< nwell >>
rect -407 -519 407 519
<< pmos >>
rect -207 -300 -177 300
rect -111 -300 -81 300
rect -15 -300 15 300
rect 81 -300 111 300
rect 177 -300 207 300
<< pdiff >>
rect -269 288 -207 300
rect -269 -288 -257 288
rect -223 -288 -207 288
rect -269 -300 -207 -288
rect -177 288 -111 300
rect -177 -288 -161 288
rect -127 -288 -111 288
rect -177 -300 -111 -288
rect -81 288 -15 300
rect -81 -288 -65 288
rect -31 -288 -15 288
rect -81 -300 -15 -288
rect 15 288 81 300
rect 15 -288 31 288
rect 65 -288 81 288
rect 15 -300 81 -288
rect 111 288 177 300
rect 111 -288 127 288
rect 161 -288 177 288
rect 111 -300 177 -288
rect 207 288 269 300
rect 207 -288 223 288
rect 257 -288 269 288
rect 207 -300 269 -288
<< pdiffc >>
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
<< nsubdiff >>
rect -371 449 -275 483
rect 275 449 371 483
rect -371 -449 -337 449
rect 337 -449 371 449
rect -371 -483 371 -449
<< nsubdiffcont >>
rect -275 449 275 483
<< poly >>
rect -129 381 -63 397
rect -129 347 -113 381
rect -79 347 -63 381
rect -129 331 -63 347
rect 63 381 129 397
rect 63 347 79 381
rect 113 347 129 381
rect 63 331 129 347
rect -207 300 -177 326
rect -111 300 -81 331
rect -15 300 15 326
rect 81 300 111 331
rect 177 300 207 326
rect -207 -331 -177 -300
rect -111 -326 -81 -300
rect -15 -331 15 -300
rect 81 -326 111 -300
rect 177 -331 207 -300
rect -225 -347 -159 -331
rect -225 -381 -209 -347
rect -175 -381 -159 -347
rect -225 -397 -159 -381
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect 159 -347 225 -331
rect 159 -381 175 -347
rect 209 -381 225 -347
rect 159 -397 225 -381
<< polycont >>
rect -113 347 -79 381
rect 79 347 113 381
rect -209 -381 -175 -347
rect -17 -381 17 -347
rect 175 -381 209 -347
<< locali >>
rect -291 449 -275 483
rect 275 449 291 483
rect -129 347 -113 381
rect -79 347 -63 381
rect 63 347 79 381
rect 113 347 129 381
rect -257 288 -223 304
rect -257 -304 -223 -288
rect -161 288 -127 304
rect -161 -304 -127 -288
rect -65 288 -31 304
rect -65 -304 -31 -288
rect 31 288 65 304
rect 31 -304 65 -288
rect 127 288 161 304
rect 127 -304 161 -288
rect 223 288 257 304
rect 223 -304 257 -288
rect -225 -381 -209 -347
rect -175 -381 -159 -347
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect 159 -381 175 -347
rect 209 -381 225 -347
<< viali >>
rect -113 347 -79 381
rect 79 347 113 381
rect -257 -288 -223 288
rect -161 -173 -127 173
rect -65 -288 -31 288
rect 31 -173 65 173
rect 127 -288 161 288
rect 223 -173 257 173
rect -209 -381 -175 -347
rect -17 -381 17 -347
rect 175 -381 209 -347
<< metal1 >>
rect -125 381 -67 387
rect 67 381 125 387
rect -125 347 -113 381
rect -79 347 79 381
rect 113 347 372 381
rect -125 341 -67 347
rect 67 341 125 347
rect -263 291 -217 300
rect -71 291 -25 300
rect 121 291 167 300
rect -263 288 167 291
rect -263 -288 -257 288
rect -223 257 -65 288
rect -223 -288 -217 257
rect -167 173 -121 185
rect -167 -134 -161 173
rect -172 -140 -161 -134
rect -127 -134 -121 173
rect -127 -140 -120 -134
rect -172 -198 -120 -192
rect -263 -300 -217 -288
rect -71 -288 -65 257
rect -31 257 127 288
rect -31 -288 -25 257
rect 25 173 71 185
rect 25 -134 31 173
rect 20 -140 31 -134
rect 65 -134 71 173
rect 65 -140 72 -134
rect 20 -198 72 -192
rect -71 -300 -25 -288
rect 121 -288 127 257
rect 161 -288 167 288
rect 217 173 263 185
rect 217 -140 223 173
rect 257 -134 263 173
rect 257 -140 270 -134
rect 212 -192 218 -140
rect 270 -192 276 -140
rect 218 -198 270 -192
rect 121 -300 167 -288
rect -221 -347 -163 -341
rect -221 -381 -209 -347
rect -175 -348 -163 -347
rect -29 -347 29 -341
rect -29 -348 -17 -347
rect -175 -381 -17 -348
rect 17 -348 29 -347
rect 163 -347 221 -341
rect 163 -348 175 -347
rect 17 -381 175 -348
rect 209 -348 221 -347
rect 338 -348 372 347
rect 209 -381 372 -348
rect -221 -382 372 -381
rect -221 -387 -163 -382
rect -29 -387 29 -382
rect 163 -387 221 -382
<< via1 >>
rect -172 -173 -161 -140
rect -161 -173 -127 -140
rect -127 -173 -120 -140
rect -172 -192 -120 -173
rect 20 -173 31 -140
rect 31 -173 65 -140
rect 65 -173 72 -140
rect 20 -192 72 -173
rect 218 -173 223 -140
rect 223 -173 257 -140
rect 257 -173 270 -140
rect 218 -192 270 -173
<< metal2 >>
rect 218 -140 270 -134
rect -178 -192 -172 -140
rect -120 -149 -114 -140
rect 14 -149 20 -140
rect -120 -183 20 -149
rect -120 -192 -114 -183
rect 14 -192 20 -183
rect 72 -149 78 -140
rect 212 -149 218 -140
rect 72 -183 218 -149
rect 72 -192 78 -183
rect 212 -192 218 -183
rect 270 -192 276 -140
rect 218 -198 270 -192
<< labels >>
flabel metal1 -258 257 160 291 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal2 s -120 -183 20 -149 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel metal1 113 347 372 381 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel nsubdiffcont 2 465 2 465 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -354 -466 354 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
