magic
tech sky130B
magscale 1 2
timestamp 1714698238
<< error_p >>
rect -29 1040 29 1046
rect -29 1006 -17 1040
rect -29 1000 29 1006
rect -125 430 -67 436
rect 67 430 125 436
rect -125 396 -113 430
rect 67 396 79 430
rect -125 390 -67 396
rect 67 390 125 396
rect -125 322 -67 328
rect 67 322 125 328
rect -125 288 -113 322
rect 67 288 79 322
rect -125 282 -67 288
rect 67 282 125 288
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect -29 -328 29 -322
rect -29 -396 29 -390
rect -29 -430 -17 -396
rect -29 -436 29 -430
rect -125 -1006 -67 -1000
rect 67 -1006 125 -1000
rect -125 -1040 -113 -1006
rect 67 -1040 79 -1006
rect -125 -1046 -67 -1040
rect 67 -1046 125 -1040
<< pwell >>
rect -311 -1178 311 1178
<< nmos >>
rect -111 468 -81 968
rect -15 468 15 968
rect 81 468 111 968
rect -111 -250 -81 250
rect -15 -250 15 250
rect 81 -250 111 250
rect -111 -968 -81 -468
rect -15 -968 15 -468
rect 81 -968 111 -468
<< ndiff >>
rect -173 956 -111 968
rect -173 480 -161 956
rect -127 480 -111 956
rect -173 468 -111 480
rect -81 956 -15 968
rect -81 480 -65 956
rect -31 480 -15 956
rect -81 468 -15 480
rect 15 956 81 968
rect 15 480 31 956
rect 65 480 81 956
rect 15 468 81 480
rect 111 956 173 968
rect 111 480 127 956
rect 161 480 173 956
rect 111 468 173 480
rect -173 238 -111 250
rect -173 -238 -161 238
rect -127 -238 -111 238
rect -173 -250 -111 -238
rect -81 238 -15 250
rect -81 -238 -65 238
rect -31 -238 -15 238
rect -81 -250 -15 -238
rect 15 238 81 250
rect 15 -238 31 238
rect 65 -238 81 238
rect 15 -250 81 -238
rect 111 238 173 250
rect 111 -238 127 238
rect 161 -238 173 238
rect 111 -250 173 -238
rect -173 -480 -111 -468
rect -173 -956 -161 -480
rect -127 -956 -111 -480
rect -173 -968 -111 -956
rect -81 -480 -15 -468
rect -81 -956 -65 -480
rect -31 -956 -15 -480
rect -81 -968 -15 -956
rect 15 -480 81 -468
rect 15 -956 31 -480
rect 65 -956 81 -480
rect 15 -968 81 -956
rect 111 -480 173 -468
rect 111 -956 127 -480
rect 161 -956 173 -480
rect 111 -968 173 -956
<< ndiffc >>
rect -161 480 -127 956
rect -65 480 -31 956
rect 31 480 65 956
rect 127 480 161 956
rect -161 -238 -127 238
rect -65 -238 -31 238
rect 31 -238 65 238
rect 127 -238 161 238
rect -161 -956 -127 -480
rect -65 -956 -31 -480
rect 31 -956 65 -480
rect 127 -956 161 -480
<< psubdiff >>
rect -275 1108 275 1142
rect -275 -1108 -241 1108
rect 241 -1108 275 1108
rect -275 -1142 -179 -1108
rect 179 -1142 275 -1108
<< psubdiffcont >>
rect -179 -1142 179 -1108
<< poly >>
rect -33 1040 33 1056
rect -33 1006 -17 1040
rect 17 1006 33 1040
rect -111 968 -81 994
rect -33 990 33 1006
rect -15 968 15 990
rect 81 968 111 994
rect -111 446 -81 468
rect -129 430 -63 446
rect -15 442 15 468
rect 81 446 111 468
rect -129 396 -113 430
rect -79 396 -63 430
rect -129 380 -63 396
rect 63 430 129 446
rect 63 396 79 430
rect 113 396 129 430
rect 63 380 129 396
rect -129 322 -63 338
rect -129 288 -113 322
rect -79 288 -63 322
rect -129 272 -63 288
rect 63 322 129 338
rect 63 288 79 322
rect 113 288 129 322
rect -111 250 -81 272
rect -15 250 15 276
rect 63 272 129 288
rect 81 250 111 272
rect -111 -276 -81 -250
rect -15 -272 15 -250
rect -33 -288 33 -272
rect 81 -276 111 -250
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -338 33 -322
rect -33 -396 33 -380
rect -33 -430 -17 -396
rect 17 -430 33 -396
rect -111 -468 -81 -442
rect -33 -446 33 -430
rect -15 -468 15 -446
rect 81 -468 111 -442
rect -111 -990 -81 -968
rect -129 -1006 -63 -990
rect -15 -994 15 -968
rect 81 -990 111 -968
rect -129 -1040 -113 -1006
rect -79 -1040 -63 -1006
rect -129 -1056 -63 -1040
rect 63 -1006 129 -990
rect 63 -1040 79 -1006
rect 113 -1040 129 -1006
rect 63 -1056 129 -1040
<< polycont >>
rect -17 1006 17 1040
rect -113 396 -79 430
rect 79 396 113 430
rect -113 288 -79 322
rect 79 288 113 322
rect -17 -322 17 -288
rect -17 -430 17 -396
rect -113 -1040 -79 -1006
rect 79 -1040 113 -1006
<< locali >>
rect -33 1006 -17 1040
rect 17 1006 33 1040
rect -161 956 -127 972
rect -161 464 -127 480
rect -65 956 -31 972
rect -65 464 -31 480
rect 31 956 65 972
rect 31 464 65 480
rect 127 956 161 972
rect 127 464 161 480
rect -129 396 -113 430
rect -79 396 -63 430
rect 63 396 79 430
rect 113 396 129 430
rect -129 288 -113 322
rect -79 288 -63 322
rect 63 288 79 322
rect 113 288 129 322
rect -161 238 -127 254
rect -161 -254 -127 -238
rect -65 238 -31 254
rect -65 -254 -31 -238
rect 31 238 65 254
rect 31 -254 65 -238
rect 127 238 161 254
rect 127 -254 161 -238
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -430 -17 -396
rect 17 -430 33 -396
rect -161 -480 -127 -464
rect -161 -972 -127 -956
rect -65 -480 -31 -464
rect -65 -972 -31 -956
rect 31 -480 65 -464
rect 31 -972 65 -956
rect 127 -480 161 -464
rect 127 -972 161 -956
rect -129 -1040 -113 -1006
rect -79 -1040 -63 -1006
rect 63 -1040 79 -1006
rect 113 -1040 129 -1006
rect -195 -1142 -179 -1108
rect 179 -1142 195 -1108
<< viali >>
rect -17 1006 17 1040
rect -161 528 -127 908
rect -65 575 -31 861
rect 31 528 65 908
rect 127 575 161 861
rect -113 396 -79 430
rect 79 396 113 430
rect -113 288 -79 322
rect 79 288 113 322
rect -161 -190 -127 190
rect -65 -143 -31 143
rect 31 -190 65 190
rect 127 -143 161 143
rect -17 -322 17 -288
rect -17 -430 17 -396
rect -161 -908 -127 -528
rect -65 -861 -31 -575
rect 31 -908 65 -528
rect 127 -861 161 -575
rect -113 -1040 -79 -1006
rect 79 -1040 113 -1006
<< metal1 >>
rect -29 1040 29 1046
rect -29 1006 -17 1040
rect 17 1006 29 1040
rect -29 1000 29 1006
rect -167 908 -121 920
rect -167 528 -161 908
rect -127 528 -121 908
rect 25 908 71 920
rect -71 861 -25 873
rect -71 575 -65 861
rect -31 575 -25 861
rect -71 563 -25 575
rect -167 516 -121 528
rect 25 528 31 908
rect 65 528 71 908
rect 121 861 167 873
rect 121 575 127 861
rect 161 575 167 861
rect 121 563 167 575
rect 25 516 71 528
rect -125 430 -67 436
rect -125 396 -113 430
rect -79 396 -67 430
rect -125 390 -67 396
rect 67 430 125 436
rect 67 396 79 430
rect 113 396 125 430
rect 67 390 125 396
rect -125 322 -67 328
rect -125 288 -113 322
rect -79 288 -67 322
rect -125 282 -67 288
rect 67 322 125 328
rect 67 288 79 322
rect 113 288 125 322
rect 67 282 125 288
rect -167 190 -121 202
rect -167 -190 -161 190
rect -127 -190 -121 190
rect 25 190 71 202
rect -71 143 -25 155
rect -71 -143 -65 143
rect -31 -143 -25 143
rect -71 -155 -25 -143
rect -167 -202 -121 -190
rect 25 -190 31 190
rect 65 -190 71 190
rect 121 143 167 155
rect 121 -143 127 143
rect 161 -143 167 143
rect 121 -155 167 -143
rect 25 -202 71 -190
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect 17 -322 29 -288
rect -29 -328 29 -322
rect -29 -396 29 -390
rect -29 -430 -17 -396
rect 17 -430 29 -396
rect -29 -436 29 -430
rect -167 -528 -121 -516
rect -167 -908 -161 -528
rect -127 -908 -121 -528
rect 25 -528 71 -516
rect -71 -575 -25 -563
rect -71 -861 -65 -575
rect -31 -861 -25 -575
rect -71 -873 -25 -861
rect -167 -920 -121 -908
rect 25 -908 31 -528
rect 65 -908 71 -528
rect 121 -575 167 -563
rect 121 -861 127 -575
rect 161 -861 167 -575
rect 121 -873 167 -861
rect 25 -920 71 -908
rect -125 -1006 -67 -1000
rect -125 -1040 -113 -1006
rect -79 -1040 -67 -1006
rect -125 -1046 -67 -1040
rect 67 -1006 125 -1000
rect 67 -1040 79 -1006
rect 113 -1040 125 -1006
rect 67 -1046 125 -1040
<< properties >>
string FIXED_BBOX -258 -1125 258 1125
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 3 nf 3 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
