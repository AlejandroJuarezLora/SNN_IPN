*MADE BY JORGE ALEJANDRO JUAREZ LORA IPN

.subckt rram_v0 TE BE
N1 TE BE rram_v0_model
.ends rram_v0

.model rram_v0_model rram_v0_va
+ g0 = 0.2751
+ V0 = 0.430 
+ I0 = 6.140e-5
+ maxGap = 1.7
+ minGap = 0.1
+ Vel0 = 150 
+ Beta0 = -1.25
+ gamma0 = 16.5
+ Ea = 0.6
+ a0 = 0.25
+ tox = 5.0
+ maxslope = 1e12
+ smoothing = 1e-8
+ GMIN = 1e-12
+ Kclip = 200


.control
pre_osdi /home/alex/pdk/sky130B/libs.tech/ngspice/rram_v0.osdi
.endc
