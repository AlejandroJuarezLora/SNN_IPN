magic
tech sky130B
magscale 1 2
timestamp 1714760917
<< error_p >>
rect -125 681 -67 687
rect 67 681 125 687
rect -125 647 -113 681
rect 67 647 79 681
rect -125 641 -67 647
rect 67 641 125 647
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -125 -647 -67 -641
rect 67 -647 125 -641
rect -125 -681 -113 -647
rect 67 -681 79 -647
rect -125 -687 -67 -681
rect 67 -687 125 -681
<< pwell >>
rect -311 -819 311 819
<< nmos >>
rect -111 109 -81 609
rect -15 109 15 609
rect 81 109 111 609
rect -111 -609 -81 -109
rect -15 -609 15 -109
rect 81 -609 111 -109
<< ndiff >>
rect -173 597 -111 609
rect -173 121 -161 597
rect -127 121 -111 597
rect -173 109 -111 121
rect -81 597 -15 609
rect -81 121 -65 597
rect -31 121 -15 597
rect -81 109 -15 121
rect 15 597 81 609
rect 15 121 31 597
rect 65 121 81 597
rect 15 109 81 121
rect 111 597 173 609
rect 111 121 127 597
rect 161 121 173 597
rect 111 109 173 121
rect -173 -121 -111 -109
rect -173 -597 -161 -121
rect -127 -597 -111 -121
rect -173 -609 -111 -597
rect -81 -121 -15 -109
rect -81 -597 -65 -121
rect -31 -597 -15 -121
rect -81 -609 -15 -597
rect 15 -121 81 -109
rect 15 -597 31 -121
rect 65 -597 81 -121
rect 15 -609 81 -597
rect 111 -121 173 -109
rect 111 -597 127 -121
rect 161 -597 173 -121
rect 111 -609 173 -597
<< ndiffc >>
rect -161 121 -127 597
rect -65 121 -31 597
rect 31 121 65 597
rect 127 121 161 597
rect -161 -597 -127 -121
rect -65 -597 -31 -121
rect 31 -597 65 -121
rect 127 -597 161 -121
<< psubdiff >>
rect -275 749 275 783
rect -275 -749 -241 749
rect 241 687 275 749
rect 241 -749 275 -687
rect -275 -783 275 -749
<< psubdiffcont >>
rect 241 -687 275 687
<< poly >>
rect -129 681 -63 697
rect -129 647 -113 681
rect -79 647 -63 681
rect -129 631 -63 647
rect 63 681 129 697
rect 63 647 79 681
rect 113 647 129 681
rect -111 609 -81 631
rect -15 609 15 635
rect 63 631 129 647
rect 81 609 111 631
rect -111 83 -81 109
rect -15 87 15 109
rect -33 71 33 87
rect 81 83 111 109
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -111 -109 -81 -83
rect -33 -87 33 -71
rect -15 -109 15 -87
rect 81 -109 111 -83
rect -111 -631 -81 -609
rect -129 -647 -63 -631
rect -15 -635 15 -609
rect 81 -631 111 -609
rect -129 -681 -113 -647
rect -79 -681 -63 -647
rect -129 -697 -63 -681
rect 63 -647 129 -631
rect 63 -681 79 -647
rect 113 -681 129 -647
rect 63 -697 129 -681
<< polycont >>
rect -113 647 -79 681
rect 79 647 113 681
rect -17 37 17 71
rect -17 -71 17 -37
rect -113 -681 -79 -647
rect 79 -681 113 -647
<< locali >>
rect 241 687 275 703
rect -129 647 -113 681
rect -79 647 -63 681
rect 63 647 79 681
rect 113 647 129 681
rect -161 597 -127 613
rect -161 105 -127 121
rect -65 597 -31 613
rect -65 105 -31 121
rect 31 597 65 613
rect 31 105 65 121
rect 127 597 161 613
rect 127 105 161 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -161 -121 -127 -105
rect -161 -613 -127 -597
rect -65 -121 -31 -105
rect -65 -613 -31 -597
rect 31 -121 65 -105
rect 31 -613 65 -597
rect 127 -121 161 -105
rect 127 -613 161 -597
rect -129 -681 -113 -647
rect -79 -681 -63 -647
rect 63 -681 79 -647
rect 113 -681 129 -647
rect 241 -703 275 -687
<< viali >>
rect -113 647 -79 681
rect 79 647 113 681
rect -161 145 -127 573
rect -65 216 -31 502
rect 31 145 65 573
rect 127 216 161 502
rect -17 37 17 71
rect -17 -71 17 -37
rect -161 -573 -127 -145
rect -65 -502 -31 -216
rect 31 -573 65 -145
rect 127 -502 161 -216
rect -113 -681 -79 -647
rect 79 -681 113 -647
<< metal1 >>
rect -125 681 -67 687
rect -125 647 -113 681
rect -79 647 -67 681
rect -125 641 -67 647
rect 67 681 125 687
rect 67 647 79 681
rect 113 647 125 681
rect 67 641 125 647
rect -167 573 -121 585
rect -167 145 -161 573
rect -127 145 -121 573
rect 25 573 71 585
rect -71 502 -25 514
rect -71 216 -65 502
rect -31 216 -25 502
rect -71 204 -25 216
rect -167 133 -121 145
rect 25 145 31 573
rect 65 145 71 573
rect 121 502 167 514
rect 121 216 127 502
rect 161 216 167 502
rect 121 204 167 216
rect 25 133 71 145
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -167 -145 -121 -133
rect -167 -573 -161 -145
rect -127 -573 -121 -145
rect 25 -145 71 -133
rect -71 -216 -25 -204
rect -71 -502 -65 -216
rect -31 -502 -25 -216
rect -71 -514 -25 -502
rect -167 -585 -121 -573
rect 25 -573 31 -145
rect 65 -573 71 -145
rect 121 -216 167 -204
rect 121 -502 127 -216
rect 161 -502 167 -216
rect 121 -514 167 -502
rect 25 -585 71 -573
rect -125 -647 -67 -641
rect -125 -681 -113 -647
rect -79 -681 -67 -647
rect -125 -687 -67 -681
rect 67 -647 125 -641
rect 67 -681 79 -647
rect 113 -681 125 -647
rect 67 -687 125 -681
<< properties >>
string FIXED_BBOX -258 -766 258 766
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 90 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
