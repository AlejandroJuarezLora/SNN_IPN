magic
tech sky130B
magscale 1 2
timestamp 1715032571
<< locali >>
rect -886 -384 271 -350
rect -1288 -1218 -1254 -1191
rect -1340 -1225 -1254 -1218
rect -1340 -1252 -1255 -1225
rect -1340 -1439 -1306 -1252
rect -886 -1439 -852 -384
rect 1158 -1253 1232 -1219
rect 744 -1439 778 -1285
rect 1198 -1439 1232 -1253
rect -1340 -1473 1232 -1439
<< viali >>
rect -21 1207 13 1241
rect -302 1075 -268 1109
rect 189 1077 223 1111
<< metal1 >>
rect -21 1253 13 1328
rect -27 1241 19 1253
rect -222 1207 -21 1241
rect 13 1240 19 1241
rect 13 1207 126 1240
rect -314 1109 -256 1115
rect -222 1109 -188 1207
rect -27 1206 126 1207
rect -27 1195 19 1206
rect -314 1075 -302 1109
rect -268 1075 -188 1109
rect -314 1069 -256 1075
rect -222 891 -188 1075
rect -21 1049 13 1195
rect 92 1111 126 1206
rect 177 1111 235 1117
rect 92 1077 189 1111
rect 223 1077 235 1111
rect 177 1071 235 1077
rect -338 857 -188 891
rect -1535 738 -1354 770
rect -102 681 -74 791
rect 1267 762 1456 798
rect -60 681 -32 685
rect -395 653 369 681
rect -60 460 -32 653
rect -882 432 772 460
rect -1438 7 -1014 42
rect -1395 -567 -1360 7
rect -882 -126 -854 432
rect -5 362 671 363
rect -779 328 671 362
rect -779 206 -745 328
rect -676 244 -154 272
rect -672 242 -438 244
rect -672 236 -440 242
rect -386 206 -334 212
rect -778 158 -745 206
rect -1000 -154 -853 -126
rect -779 -249 -745 158
rect -590 154 -584 206
rect -532 154 -526 206
rect -386 148 -334 154
rect -186 100 -158 244
rect 18 232 24 284
rect 76 272 82 284
rect 76 266 270 272
rect 76 244 466 266
rect 76 232 82 244
rect 230 236 466 244
rect 528 207 580 213
rect 307 155 313 207
rect 365 155 371 207
rect 528 149 580 155
rect -187 48 -156 100
rect -187 17 -39 48
rect -186 -98 -158 17
rect -186 -126 66 -98
rect -89 -241 -83 -229
rect -779 -283 -391 -249
rect -182 -269 -83 -241
rect -1011 -478 -1005 -466
rect -1294 -506 -1005 -478
rect -1011 -518 -1005 -506
rect -953 -518 -947 -466
rect -1395 -602 -1106 -567
rect -781 -591 -295 -557
rect -1395 -1484 -1360 -602
rect -1147 -713 -847 -675
rect -1201 -843 -1149 -837
rect -1005 -843 -953 -837
rect -1011 -895 -1005 -843
rect -953 -895 -947 -843
rect -1201 -901 -1149 -895
rect -1005 -901 -953 -895
rect -1291 -1224 -1061 -1196
rect -1240 -1322 -1008 -1284
rect -1240 -1389 -1202 -1322
rect -885 -1389 -847 -713
rect -781 -1289 -747 -591
rect -182 -666 -154 -269
rect -89 -281 -83 -269
rect -31 -281 -25 -229
rect 38 -666 66 -126
rect 636 -248 670 328
rect 744 -126 772 432
rect 1257 43 1295 45
rect 888 5 1327 43
rect 742 -158 897 -126
rect 282 -282 670 -248
rect 636 -559 670 -282
rect 839 -522 845 -470
rect 897 -482 903 -470
rect 897 -510 1176 -482
rect 897 -522 903 -510
rect 185 -593 670 -559
rect -671 -692 -154 -666
rect -671 -696 -170 -692
rect 28 -696 466 -666
rect -579 -896 -527 -890
rect -387 -896 -335 -890
rect -192 -896 -140 -890
rect 128 -892 180 -886
rect -393 -948 -387 -896
rect -335 -948 -329 -896
rect -198 -948 -192 -896
rect -140 -948 -134 -896
rect -579 -954 -527 -948
rect -387 -954 -335 -948
rect -192 -954 -140 -948
rect 128 -950 180 -944
rect 325 -892 377 -886
rect 325 -950 377 -944
rect 513 -892 565 -886
rect 513 -950 565 -944
rect 636 -1289 670 -593
rect -781 -1323 670 -1289
rect 738 -567 776 -563
rect 1257 -567 1295 5
rect 738 -605 1295 -567
rect 738 -1389 776 -605
rect 995 -712 1288 -676
rect 1040 -857 1092 -851
rect 839 -909 845 -857
rect 897 -909 903 -857
rect 1040 -915 1092 -909
rect 953 -1225 1181 -1192
rect 1251 -1285 1288 -712
rect 903 -1322 1288 -1285
rect -1240 -1427 776 -1389
rect 1251 -1484 1288 -1322
rect -1395 -1519 1289 -1484
rect -1395 -1523 -1360 -1519
rect 1251 -1520 1288 -1519
<< via1 >>
rect -584 154 -532 206
rect -386 154 -334 206
rect 24 232 76 284
rect 313 155 365 207
rect 528 155 580 207
rect -1005 -518 -953 -466
rect -1201 -895 -1149 -843
rect -1005 -895 -953 -843
rect -83 -281 -31 -229
rect 845 -522 897 -470
rect -579 -948 -527 -896
rect -387 -948 -335 -896
rect -192 -948 -140 -896
rect 128 -944 180 -892
rect 325 -944 377 -892
rect 513 -944 565 -892
rect 845 -909 897 -857
rect 1040 -909 1092 -857
<< metal2 >>
rect 24 284 76 290
rect 24 226 76 232
rect -584 206 -532 212
rect -778 166 -584 194
rect -778 -370 -750 166
rect -392 194 -386 206
rect -532 166 -386 194
rect -392 154 -386 166
rect -334 154 -328 206
rect 35 195 64 226
rect 313 207 365 213
rect -584 148 -532 154
rect 35 48 63 195
rect 522 196 528 207
rect 365 166 528 196
rect 522 155 528 166
rect 580 196 586 207
rect 580 166 667 196
rect 580 155 586 166
rect 313 149 365 155
rect -71 20 63 48
rect -83 -229 -31 -223
rect 35 -241 63 20
rect -31 -269 63 -241
rect -83 -287 -31 -281
rect -860 -398 -750 -370
rect 637 -398 667 166
rect -1005 -466 -953 -460
rect -1005 -524 -953 -518
rect -993 -624 -965 -524
rect -860 -624 -832 -398
rect -993 -652 -832 -624
rect -993 -837 -965 -652
rect -1005 -843 -953 -837
rect -1207 -895 -1201 -843
rect -1149 -855 -1143 -843
rect -1011 -855 -1005 -843
rect -1149 -883 -1005 -855
rect -1149 -895 -1143 -883
rect -1011 -895 -1005 -883
rect -953 -895 -947 -843
rect -1005 -901 -953 -895
rect -778 -908 -750 -398
rect 636 -426 741 -398
rect 637 -427 741 -426
rect -387 -896 -335 -890
rect -192 -896 -140 -890
rect -585 -908 -579 -896
rect -782 -936 -579 -908
rect -585 -948 -579 -936
rect -527 -908 -521 -896
rect -393 -908 -387 -896
rect -527 -936 -387 -908
rect -527 -948 -521 -936
rect -393 -948 -387 -936
rect -335 -908 -329 -896
rect -198 -908 -192 -896
rect -335 -936 -192 -908
rect -335 -948 -329 -936
rect -198 -948 -192 -936
rect -140 -948 -134 -896
rect 122 -944 128 -892
rect 180 -903 186 -892
rect 319 -903 325 -892
rect 180 -933 325 -903
rect 180 -944 186 -933
rect 319 -944 325 -933
rect 377 -903 383 -892
rect 507 -903 513 -892
rect 377 -933 513 -903
rect 377 -944 383 -933
rect 507 -944 513 -933
rect 565 -903 571 -892
rect 637 -903 667 -427
rect 713 -620 741 -427
rect 845 -470 897 -464
rect 845 -528 897 -522
rect 857 -620 885 -528
rect 713 -648 885 -620
rect 857 -851 885 -648
rect 565 -933 667 -903
rect 845 -857 897 -851
rect 1034 -869 1040 -857
rect 897 -897 1040 -869
rect 1034 -909 1040 -897
rect 1092 -909 1098 -857
rect 845 -915 897 -909
rect 565 -944 571 -933
rect -387 -954 -335 -948
rect -192 -954 -140 -948
use rram2_0  rram2_0_0
timestamp 1714756818
transform 1 0 -58 0 1 32
box -32 -32 32 32
use sky130_fd_pr__nfet_01v8_AKC4V5  sky130_fd_pr__nfet_01v8_AKC4V5_0
timestamp 1714760917
transform -1 0 1017 0 1 -639
box -311 -819 311 819
use sky130_fd_pr__nfet_01v8_AKC4V5  sky130_fd_pr__nfet_01v8_AKC4V5_1
timestamp 1714760917
transform 1 0 -1127 0 1 -639
box -311 -819 311 819
use sky130_fd_pr__nfet_01v8_JZLRWN  sky130_fd_pr__nfet_01v8_JZLRWN_0
timestamp 1714757534
transform 1 0 395 0 1 40
box -311 -460 311 460
use sky130_fd_pr__nfet_01v8_JZLRWN  sky130_fd_pr__nfet_01v8_JZLRWN_1
timestamp 1714757534
transform 1 0 -505 0 1 40
box -311 -460 311 460
use sky130_fd_pr__pfet_01v8_86T979  sky130_fd_pr__pfet_01v8_86T979_0
timestamp 1715032421
transform 1 0 -48 0 1 893
box -211 -384 211 384
use sky130_fd_pr__pfet_01v8_R4E532  sky130_fd_pr__pfet_01v8_R4E532_0
timestamp 1714756698
transform 1 0 299 0 1 -939
box -407 -519 407 519
use sky130_fd_pr__pfet_01v8_R4E532  sky130_fd_pr__pfet_01v8_R4E532_1
timestamp 1714756698
transform 1 0 -409 0 1 -939
box -407 -519 407 519
use sky130_fd_pr__pfet_01v8_RWS95J  sky130_fd_pr__pfet_01v8_RWS95J_0
timestamp 1714698450
transform 1 0 -845 0 1 828
box -696 -319 696 319
use sky130_fd_pr__pfet_01v8_RWS95J  sky130_fd_pr__pfet_01v8_RWS95J_1
timestamp 1714698450
transform 1 0 761 0 1 826
box -696 -319 696 319
<< labels >>
flabel metal1 s -137 29 -137 29 0 FreeSans 640 0 0 0 BE
flabel metal2 s 42 34 42 34 0 FreeSans 640 0 0 0 TE
flabel metal2 s -866 -411 -838 -383 0 FreeSans 640 0 0 0 vpre
flabel metal2 s 637 -427 745 -397 0 FreeSans 640 0 0 0 vpost
flabel metal1 s -57 346 -57 346 0 FreeSans 640 0 0 0 R
flabel metal1 s 1311 23 1311 23 0 FreeSans 640 0 0 0 vout_post
port 1 nsew
flabel metal1 s -1438 7 -1403 42 0 FreeSans 640 0 0 0 vout_pre
port 2 nsew
flabel locali -55 -1456 -55 -1456 0 FreeSans 640 0 0 0 gnd
port 3 nsew
flabel metal1 -51 447 -51 447 0 FreeSans 640 0 0 0 Im10
flabel metal1 -5 1300 -5 1300 0 FreeSans 640 0 0 0 VDD
port 4 nsew
flabel metal1 -1517 753 -1517 753 0 FreeSans 640 0 0 0 I_pre
port 5 nsew
flabel metal1 1431 781 1431 781 0 FreeSans 640 0 0 0 I_post
port 6 nsew
<< end >>
