** sch_path: /home/alex/Desktop/EDA/SNN_IPN/tb_4x8x4.sch
**.subckt tb_4x8x4
Vdd VDD GND 1.8
x1 VDD GND x N1 N2 N3 N4 layer_input
x2 VDD net10 GND net11 net12 net1 net13 M1 M2 M3 M4 layer_output
x3 VDD net15 hx x Vr1 GND opamp_sky130
R2 hx GND 9k m=1
I0 net15 GND 100u
Vin1 x net16 SINE(0 0.3 200 0 0 0)
Vread net1 net2 0
Vin3 net16 net17 SINE(0 0.5 500 0 0 90)
Vin4 net17 GND 0.9
x4 VDD net9 GND net8 net7 J1 J2 net6 J3 net5 J4 net4 J5 net3 J6 J7 net14 J8 layer_hidden
x5 VDD net9 net8 net7 GND J1 J2 net3 net14 net5 J3 net6 net4 J8 J7 J6 J5 J4 N1 N2 N3 N4 stdp_4x8
x6 Vr1 net11 net10 M2 net12 GND M1 M3 net13 M4 J1 J2 J3 J4 J5 J6 J7 J8 VDD rstdp_array_8x4
R1 net2 hx 9k m=1
**** begin user architecture code

** opencircuitdesign pdks install
.inc ~/pdk/sky130B/libs.tech/ngspice/rram_v0.spice
**.inc ~/pdk/sky130B/libs.tech/ngspice/sky.spice



.param mc_mm_switch=0
.param mc_pr_switch=0
.include ~/pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include ~/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice


**** end user architecture code
**.ends

* expanding   symbol:  layer/layer_input.sym # of pins=7
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_input.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_input.sch
.subckt layer_input vdd vss vin vout1 vout2 vout3 vout4
*.iopin vdd
*.iopin vss
*.ipin vin
*.iopin vout1
*.iopin vout2
*.iopin vout3
*.iopin vout4
x6 net2 vdd vg100n vout1 net1 vss ul_tun
x4 vdd vin net6 vss syn_pos
x8 vdd vin net2 vss syn_neg
I9 vg100n vss 100nA
XM4 vg100n vg100n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vileak vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I1 vdd vileak 100nA
x1 net4 vdd vg100n vout2 net3 vss ul_tun
x2 vdd vin net4 vss syn_neg
XM3 net3 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x3 net6 vdd vg100n vout3 net5 vss ul_tun
XM5 net5 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x7 vdd vin net8 vss syn_pos
x9 net8 vdd vg100n vout4 net7 vss ul_tun
XM6 net7 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  layer/layer_output.sym # of pins=11
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_output.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_output.sch
.subckt layer_output vdd Iext1 vss Iext2 Iext3 Iout Iext4 vout1 vout2 vout3 vout4
*.iopin vdd
*.iopin vss
*.ipin Iext1
*.iopin Iout
*.ipin Iext2
*.ipin Iext3
*.ipin Iext4
*.iopin vout1
*.iopin vout2
*.iopin vout3
*.iopin vout4
x6 Iext1 vdd vg100n vout1 net1 vss ul_tun
I9 vg100n vss 100nA
XM4 vg100n vg100n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vileak vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I1 vdd vileak 100nA
x1 Iext2 vdd vg100n vout2 net2 vss ul_tun
XM3 net2 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x3 Iext3 vdd vg100n vout3 net3 vss ul_tun
XM5 net3 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x9 Iext4 vdd vg100n vout4 net4 vss ul_tun
XM6 net4 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x14 VDD Iout net5 GND integrator
XM7 net5 vout1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net5 vout2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net5 vout3 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net5 vout4 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  OPAMP/opamp_sky130.sym # of pins=6
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/OPAMP/opamp_sky130.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/OPAMP/opamp_sky130.sch
.subckt opamp_sky130 vdd iref vin_n vin_p vout vss
*.iopin vdd
*.iopin vss
*.ipin vin_n
*.ipin vin_p
*.ipin iref
*.opin vout
XM1 vbn vin_n vp vp sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=200 m=200
XM2 voe1 vin_p vp vp sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=200 m=200
XM3 vbn vbn vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=30 m=30
XM4 voe1 vbn vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=30 m=30
XM5 vp iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=30 m=30
XM7 vout iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=150 m=150
XM8 iref iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=15 m=15
XM9 net1 vdd voe1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
XC1 net1 vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 MF=6 m=6
XM6 vout voe1 vss vss sky130_fd_pr__nfet_01v8 L=0.45 W=4.5 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=150 m=150
.ends


* expanding   symbol:  layer/layer_hidden.sym # of pins=18
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_hidden.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/layer/layer_hidden.sch
.subckt layer_hidden vdd Iext1 vss Iext2 Iext3 vout1 vout2 Iext4 vout3 Iext5 vout4 Iext6 vout5 Iext7 vout6 vout7 Iext8 vout8
*.iopin vdd
*.iopin vss
*.ipin Iext1
*.ipin Iext2
*.ipin Iext3
*.ipin Iext4
*.iopin vout1
*.iopin vout2
*.iopin vout3
*.iopin vout4
*.ipin Iext5
*.ipin Iext6
*.ipin Iext7
*.iopin Iext8
*.iopin vout5
*.iopin vout6
*.iopin vout7
*.iopin vout8
x6 Iext1 vdd vg100n vout1 net1 vss ul_tun
I9 vg100n vss 100nA
XM4 vg100n vg100n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vileak vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I1 vdd vileak 100nA
x1 Iext2 vdd vg100n vout2 net2 vss ul_tun
XM3 net2 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 Iext3 vdd vg100n vout3 net3 vss ul_tun
XM7 net3 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x3 Iext4 vdd vg100n vout4 net4 vss ul_tun
XM5 net4 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x4 Iext5 vdd vg100n vout5 net5 vss ul_tun
XM6 net5 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x5 Iext6 vdd vg100n vout6 net6 vss ul_tun
XM8 net6 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x7 Iext7 vdd vg100n vout7 net7 vss ul_tun
XM9 net7 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x8 Iext8 vdd vg100n vout8 net8 vss ul_tun
XM10 net8 vileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  Synapse/stdp_4x8.sym # of pins=22
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/stdp_4x8.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/stdp_4x8.sch
.subckt stdp_4x8 vdda i_post1 i_post2 i_post3 vssa vout_post1 vout_post2 i_post7 i_post8 i_post5 vout_post3 i_post4 i_post6
+ vout_post8 vout_post7 vout_post6 vout_post5 vout_post4 vout_pre1 vout_pre2 vout_pre3 vout_pre4
*.ipin vout_pre1
*.opin vout_post1
*.iopin vdda
*.iopin vssa
*.iopin i_post1
*.iopin i_post3
*.iopin i_post4
*.ipin vout_pre2
*.ipin vout_pre3
*.ipin vout_pre4
*.opin vout_post2
*.opin vout_post3
*.opin vout_post4
*.iopin i_post2
*.iopin i_post5
*.opin vout_post5
*.iopin i_post6
*.opin vout_post6
*.iopin i_post7
*.opin vout_post7
*.iopin i_post8
*.opin vout_post8
xstdp1 vdda vssa vout_pre1 vout_post1 i_post1 stdp
xstdp2 vdda vssa vout_pre1 vout_post2 i_post2 stdp
xstdp3 vdda vssa vout_pre1 vout_post3 i_post3 stdp
xstdp4 vdda vssa vout_pre1 vout_post4 i_post4 stdp
xstdp5 vdda vssa vout_pre2 vout_post1 i_post1 stdp
xstdp6 vdda vssa vout_pre2 vout_post2 i_post2 stdp
xstdp7 vdda vssa vout_pre2 vout_post3 i_post3 stdp
xstdp8 vdda vssa vout_pre2 vout_post4 i_post4 stdp
xstdp9 vdda vssa vout_pre3 vout_post1 i_post1 stdp
xstdp10 vdda vssa vout_pre3 vout_post2 i_post2 stdp
xstdp11 vdda vssa vout_pre3 vout_post3 i_post3 stdp
xstdp12 vdda vssa vout_pre3 vout_post4 i_post4 stdp
xstdp13 vdda vssa vout_pre4 vout_post1 i_post1 stdp
xstdp14 vdda vssa vout_pre4 vout_post2 i_post2 stdp
xstdp15 vdda vssa vout_pre4 vout_post3 i_post3 stdp
xstdp16 vdda vssa vout_pre4 vout_post4 i_post4 stdp
xstdp17 vdda vssa vout_pre1 vout_post5 i_post5 stdp
xstdp18 vdda vssa vout_pre1 vout_post6 i_post6 stdp
xstdp19 vdda vssa vout_pre1 vout_post7 i_post7 stdp
xstdp20 vdda vssa vout_pre1 vout_post8 i_post8 stdp
xstdp21 vdda vssa vout_pre2 vout_post5 i_post5 stdp
xstdp22 vdda vssa vout_pre2 vout_post6 i_post6 stdp
xstdp23 vdda vssa vout_pre2 vout_post7 i_post7 stdp
xstdp24 vdda vssa vout_pre2 vout_post8 i_post8 stdp
xstdp25 vdda vssa vout_pre3 vout_post5 i_post5 stdp
xstdp26 vdda vssa vout_pre3 vout_post6 i_post6 stdp
xstdp27 vdda vssa vout_pre3 vout_post7 i_post7 stdp
xstdp28 vdda vssa vout_pre3 vout_post8 i_post8 stdp
xstdp29 vdda vssa vout_pre4 vout_post5 i_post5 stdp
xstdp30 vdda vssa vout_pre4 vout_post6 i_post6 stdp
xstdp31 vdda vssa vout_pre4 vout_post7 i_post7 stdp
xstdp32 vdda vssa vout_pre4 vout_post8 i_post8 stdp
.ends


* expanding   symbol:  Synapse/rstdp_array_8x4.sym # of pins=19
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/rstdp_array_8x4.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/rstdp_array_8x4.sch
.subckt rstdp_array_8x4 Vr i_post2 i_post1 vout_post2 i_post3 vssa vout_post1 vout_post3 i_post4 vout_post4 vout_pre1 vout_pre2
+ vout_pre3 vout_pre4 vout_pre5 vout_pre6 vout_pre7 vout_pre8 vdda
*.ipin vout_pre1
*.opin vout_post1
*.iopin vdda
*.iopin vssa
*.iopin i_post1
*.iopin i_post3
*.iopin i_post4
*.ipin vout_pre2
*.ipin vout_pre3
*.ipin vout_pre4
*.opin vout_post2
*.opin vout_post3
*.opin vout_post4
*.iopin i_post2
*.iopin Vr
*.ipin vout_pre5
*.ipin vout_pre6
*.ipin vout_pre7
*.ipin vout_pre8
xrstdp1 vdda Vr vssa vout_pre1 vout_post1 i_post1 rstdp_mirror
xrstdp2 vdda Vr vssa vout_pre1 vout_post2 i_post2 rstdp_mirror
xrstdp3 vdda Vr vssa vout_pre1 vout_post3 i_post3 rstdp_mirror
xrstdp4 vdda Vr vssa vout_pre1 vout_post4 i_post4 rstdp_mirror
xrstdp5 vdda Vr vssa vout_pre2 vout_post1 i_post1 rstdp_mirror
xrstdp6 vdda Vr vssa vout_pre2 vout_post2 i_post2 rstdp_mirror
xrstdp7 vdda Vr vssa vout_pre2 vout_post3 i_post3 rstdp_mirror
xrstdp8 vdda Vr vssa vout_pre2 vout_post4 i_post4 rstdp_mirror
xrstdp9 vdda Vr vssa vout_pre3 vout_post1 i_post1 rstdp_mirror
xrstdp10 vdda Vr vssa vout_pre3 vout_post2 i_post2 rstdp_mirror
xrstdp11 vdda Vr vssa vout_pre3 vout_post3 i_post3 rstdp_mirror
xrstdp12 vdda Vr vssa vout_pre3 vout_post4 i_post4 rstdp_mirror
xrstdp13 vdda Vr vssa vout_pre4 vout_post1 i_post1 rstdp_mirror
xrstdp14 vdda Vr vssa vout_pre4 vout_post2 i_post2 rstdp_mirror
xrstdp15 vdda Vr vssa vout_pre4 vout_post3 i_post3 rstdp_mirror
xrstdp16 vdda Vr vssa vout_pre4 vout_post4 i_post4 rstdp_mirror
xrstdp17 vdda Vr vssa vout_pre5 vout_post1 i_post1 rstdp_mirror
xrstdp18 vdda Vr vssa vout_pre5 vout_post2 i_post2 rstdp_mirror
xrstdp19 vdda Vr vssa vout_pre5 vout_post3 i_post3 rstdp_mirror
xrstdp20 vdda Vr vssa vout_pre5 vout_post4 i_post4 rstdp_mirror
xrstdp21 vdda Vr vssa vout_pre6 vout_post1 i_post1 rstdp_mirror
xrstdp22 vdda Vr vssa vout_pre6 vout_post2 i_post2 rstdp_mirror
xrstdp23 vdda Vr vssa vout_pre6 vout_post3 i_post3 rstdp_mirror
xrstdp24 vdda Vr vssa vout_pre6 vout_post4 i_post4 rstdp_mirror
xrstdp25 vdda Vr vssa vout_pre7 vout_post1 i_post1 rstdp_mirror
xrstdp26 vdda Vr vssa vout_pre7 vout_post2 i_post2 rstdp_mirror
xrstdp27 vdda Vr vssa vout_pre7 vout_post3 i_post3 rstdp_mirror
xrstdp28 vdda Vr vssa vout_pre7 vout_post4 i_post4 rstdp_mirror
xrstdp29 vdda Vr vssa vout_pre8 vout_post1 i_post1 rstdp_mirror
xrstdp30 vdda Vr vssa vout_pre8 vout_post2 i_post2 rstdp_mirror
xrstdp31 vdda Vr vssa vout_pre8 vout_post3 i_post3 rstdp_mirror
xrstdp32 vdda Vr vssa vout_pre8 vout_post4 i_post4 rstdp_mirror
.ends


* expanding   symbol:  Neuron/ultralif/ul_tun.sym # of pins=6
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/ul_tun.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/ul_tun.sch
.subckt ul_tun Iext vdd g100n vout Ileak vss
*.iopin Iext
*.iopin vout
*.iopin vss
*.iopin Ileak
*.iopin vdd
*.iopin g100n
XM1 Ileak Ileak net1 vdd sky130_fd_pr__pfet_01v8 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Ileak net2 net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 Ileak vss vss sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C1 net1 vss 1p m=1
XM5 vout_n Ileak vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 vout_n g100n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 vout vout_n vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 vout vout_n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 vout Iext vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  Neuron/ultralif/syn_pos.sym # of pins=4
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/syn_pos.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/syn_pos.sch
.subckt syn_pos vdd Vin Isyn vss
*.iopin Vin
*.iopin vdd
*.iopin vss
*.iopin Isyn
XM9 Isyn vx vdd vdd sky130_fd_pr__pfet_01v8 L=1.1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 vx vx vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM12 vx Vin vss vss sky130_fd_pr__nfet_01v8 L=1 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Isyn net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net1 vdd sky130_fd_pr__res_generic_po W=1.15 L=1 m=1
R2 vss net1 sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends


* expanding   symbol:  Neuron/ultralif/syn_neg.sym # of pins=4
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/syn_neg.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/syn_neg.sch
.subckt syn_neg vdd Vin Isyn vss
*.iopin Vin
*.iopin Isyn
*.iopin vdd
*.iopin vss
XM10 Isyn Vin vx vdd sky130_fd_pr__pfet_01v8 L=35 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vx Vin vdd vdd sky130_fd_pr__pfet_01v8 L=35 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Isyn net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 net1 vdd sky130_fd_pr__res_generic_po W=1.15 L=1 m=1
R2 vss net1 sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends


* expanding   symbol:  Neuron/ultralif/integrator.sym # of pins=4
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/integrator.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Neuron/ultralif/integrator.sch
.subckt integrator vdd Iout Ispks gnd
*.iopin Ispks
*.iopin Iout
*.iopin vdd
*.iopin gnd
XMIn Ispks vx vsyn vdd sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vsyn vdd vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=24.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Iout vsyn vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=24.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XCsyn vdd vsyn sky130_fd_pr__cap_mim_m3_1 W=22.5 L=22 MF=1 m=1
R2 vx vdd sky130_fd_pr__res_generic_po W=1 L=1 m=1
R1 gnd vx sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends


* expanding   symbol:  Synapse/stdp.sym # of pins=5
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/stdp.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/stdp.sch
.subckt stdp vdd vss vout_pre vout_post I_post
*.iopin vdd
*.iopin vss
*.iopin vout_post
*.iopin vout_pre
*.iopin I_post
XM2 A vout_pre te vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 te vout_post vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 A vout_post net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 vout_pre vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR2 te be rram_v0
XM14 I_post A vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 A A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmr be net1 0
.save i(vmr)
**** begin user architecture code


.save v(te,be)


**** end user architecture code
.ends


* expanding   symbol:  Synapse/rstdp_mirror.sym # of pins=6
** sym_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/rstdp_mirror.sym
** sch_path: /home/alex/Desktop/EDA/SNN_IPN/Synapse/rstdp_mirror.sch
.subckt rstdp_mirror vdd R vss vout_pre vout_post I_post
*.iopin vdd
*.iopin vss
*.iopin R
*.iopin vout_post
*.iopin vout_pre
*.iopin I_post
XM2 A vout_pre vpre vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vpre vout_post vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 A vout_post vpost vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vpost vout_pre vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR2 be te rram_v0
XM5 vpre R te vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 R vpost vss sky130_fd_pr__nfet_01v8 L=0.15 W=7.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 vpre R net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 te R vpost vdd sky130_fd_pr__pfet_01v8 L=0.15 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 I_post A vdd vdd sky130_fd_pr__pfet_01v8 L=3 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 A A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmr be net1 0
.save i(vmr)
**** begin user architecture code


.save v(te,be)


**** end user architecture code
.ends

.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code



.options method gear
.options KLU
.options noinit
.options set num_threads=10
.options set ng_nomodcheck
.options set skywaterpdk
.options set wr_vecnames
.options set wr_singlescale
.options numdgt = 2
.save x Vr1 I(Vread) hx x
+N1 N2 N3 N4 M1 M2 M3 M4
+J1 J2 J3 J4 J5 J6 J7 J8

.tran 5u 25m 0 100n



**** end user architecture code
.end
