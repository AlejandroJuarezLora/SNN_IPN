*si le pones el valor de g0 a gap0, hay lissajous
.subckt rram_v0 TE BE PARAMS:
+Gap_0=unif(0.9,0.8)
*+Gap_0=unif(0.9,0.8)
+g0=0.2751
+V0=0.430
+I0=6.140e-5
+maxGap=1.7
+minGap=0.1
+Vel0=150
+Beta0=-1.25 
+gamma0=16.5
+Ea=1.500 
+a0=0.25
+tox=5.0 
+smoothing=1e-8
+Kclip=50
+vt=0.0258
+maxslope=1e18
+GMIN = 1e-12

* Auxiliary resistor for stable conductance
Raux r 0 1e12

* Capacitor with initial condition
Cr r 0 1 IC={Gap_0}

* Variable conductance resistor
Gr 0 r value={ddt(-1e-9 * V(r) - V(BE)) + ddt_Gap(V(TE) - V(BE),V(r)) + clip_minGap(V(r), ddt_Gap(V(TE) - V(BE), V(r))) + clip_maxGap(V(r), ddt_Gap(V(TE) - V(BE), V(r)))}

* Memristor conductance
Gpm TE BE value={I0 * safeexp(-(V(r))/g0) * safesinh((V(TE) - V(BE))/V0) }

* Function for smooth step approximation
.func smth_stp(x)={0.5*(x/sqrt(x*x + smoothing)+1)}

* Gamma function dependent on voltage
.func gamma(Gap)={gamma0+Beta0*pow(Gap,3)}

* Rate of change of gap
.func ddt_Gap(vtb, Gap)={-(maxGap - minGap) * Vel0 * safeexp(-Ea/vt) * safesinh(vtb * gamma(Gap) * a0/(tox * vt))}

* Clipping function for minimum gap
.func clip_minGap(gap, ddtGap)={(safeexp(Kclip*(minGap - gap)) - ddtGap) * smth_stp(minGap - gap)}

* Clipping function for maximum gap
.func clip_maxGap(gap, ddtGap)={(-safeexp(Kclip*(gap - maxGap)) - ddtGap) * smth_stp(gap - maxGap)}
.func safeexp(x)={exp(x*(x <= log(maxslope)))*(x <= log(maxslope)) + (x>log(maxslope))*(maxslope + maxslope*(x-log(maxslope)))}
.func safesinh(x)={0.5*(safeexp(x) - safeexp(-x))}


.ends rram_v0